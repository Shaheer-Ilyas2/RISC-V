`timescale 1ns / 1ps

module mux_4x1(
        input  logic [31:0] in1, in2, in3, in4,
        input  logic [1:0]  sel,
        output logic [31:0] out
    );
    
    always_comb begin
        if      (sel == 2'b00) out = in1;
        else if (sel == 2'b01) out = in2;
        else if (sel == 2'b10) out = in3;
        else if (sel == 2'b11) out = in4;
    end
    
endmodule